library verilog;
use verilog.vl_types.all;
entity mydisp_vlg_vec_tst is
end mydisp_vlg_vec_tst;
